-- Elementos de Sistemas
-- by Luciano Soares
-- Mux8Way.vhd

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Mux8Way is
	port ( 
			a:   in  STD_LOGIC;
			b:   in  STD_LOGIC;
			c:   in  STD_LOGIC;
			d:   in  STD_LOGIC;
			e:   in  STD_LOGIC;
			f:   in  STD_LOGIC;
			g:   in  STD_LOGIC;
			h:   in  STD_LOGIC;
			sel: in  STD_LOGIC_VECTOR(2 downto 0);
			q:   out STD_LOGIC);
end entity;

architecture arch of Mux8Way is
begin

	with sel select
	q<= a when "000",
        b when "001",
        c when "010",
        d when "011",
        e when "100",
        f when "101",
        g when "110",
        h when others;
        
end architecture;