library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BarrelShifter8 is
	port ( 
			a:   in  STD_LOGIC_VECTOR(7 downto 0);
			q:   out STD_LOGIC_VECTOR(7 downto 0));
end entity;

architecture arch of BarrelShifter8 is
begin

end main;